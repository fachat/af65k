----------------------------------------------------------------------------------
--
--    Opcode map for the af65k CPU
--
--    Copyright (C) 2011,2012 André Fachat
--
--    This library is free software; you can redistribute it and/or
--    modify it under the terms of the GNU Lesser General Public
--    License as published by the Free Software Foundation; either
--    version 2.1 of the License, or (at your option) any later version.
--
--    This library is distributed in the hope that it will be useful,
--    but WITHOUT ANY WARRANTY; without even the implied warranty of
--    MERCHANTABILITY or FITNESS FOR A PARTICULAR PURPOSE.  See the GNU
--    Lesser General Public License for more details.
--
--    You should have received a copy of the GNU Lesser General Public
--    License along with this library; if not, write to the Free Software
--    Foundation, Inc., 51 Franklin Street, Fifth Floor, Boston, MA  02110-1301  USA
--
----------------------------------------------------------------------------------
--
-- 	entity: 		af65002opmap
--		purpose:		maps bytes read into operations and addressing modes
--		features:	- main case switch is generated from an XML file (see further documentation)
--		version:		0.1 (first public release)
--		date:			18mar2012
--		
--		Changes:		
--

library IEEE;
use IEEE.STD_LOGIC_1164.ALL;
library af65002;
use af65002.af65k.all;

-- Uncomment the following library declaration if using
-- arithmetic functions with Signed or Unsigned values
--use IEEE.NUMERIC_STD.ALL;

-- Uncomment the following library declaration if instantiating
-- any Xilinx primitives in this code.
--library UNISIM;
--use UNISIM.VComponents.all;

entity af65002opmap is
   Port ( 
			opcode : in  STD_LOGIC_VECTOR (7 downto 0);
			opmap : in  STD_LOGIC_VECTOR (7 downto 0);
			prefix_rs : in rs_width;
			prefix_am : in std_logic;

			-- true when valid
			is_valid : out std_logic;
			operation : out cpu_operation;
			
			-- parameter length and syntax together define the addressing mode
			-- e.g. syntax=ABSOLUTE and adwidth=wBYTE is zeropage addressing
			-- also indwidth defines the address width for indirect addresses (only 
			-- word, long or quad
			parwidth : out par_width;
			indwidth : out rs_width;
			admode : out cpu_syntax;
			idxreg : out idx_register;
			default_le : out ext_type
	);
end af65002opmap;

architecture Behavioral of af65002opmap is

	-- opcode page
	-- 00 = std
	-- 01 = EXT
	-- 10 = QUICK
	-- 11 = SYS
	signal mapin : std_logic_vector (9 downto 0);
	
	signal pw_rs : par_width;
	signal pw_bl : par_width;
	signal pw_wq : par_width;
	
begin

	-- prepared signals
	pw_rs <= rs_width_par_width(prefix_rs);	
	pw_bl <= pBYTE when (prefix_am = '0') else pLONG;
	pw_wq <= pWORD when (prefix_am = '0') else pQUAD;

	-- input map
	mapin(9 downto 8) <= opmap(1 downto 0);
	mapin(7 downto 0) <= opcode(7 downto 0);
	
	-- generated decoding from af65002.xml
	map_p : process (mapin, pw_bl, pw_rs, pw_wq)
	begin

		operation <= xUNKNOWN;
		admode <= sUNKNOWN;
		idxreg <= iXR;			-- don't care
		indwidth <= wWORD;
		parwidth <= pNONE;
		default_le <= eNONE;
		is_valid <= '1';


case mapin is
when "0000000000" =>          -- $00, BRK Immediate: #byte 
  operation <= xBRK;
  parwidth <= pw_rs;
  admode <= sIMMEDIATE;
when "0000000001" =>          -- $01, ORA Zeropage indexed with X indirect 16bit: (zp,X) 
  operation <= xORA;
  idxreg <= iXR;
  indwidth <= wWORD;
  parwidth <= pBYTE;
  admode <= sPREINDIRECT;
when "0000000010" =>          -- $02, LDA Zeropage indexed with Y: zp,Y  (65k)
  operation <= xLDA;
  default_le <= eZERO;
  idxreg <= iYR;
  parwidth <= pw_bl;
  admode <= sABSOLUTEIND;
when "0000000011" =>          -- $03, ORA Zeropage indexed with X indirect 64bit: [[zp,X]]  (65k)
  operation <= xORA;
  idxreg <= iXR;
  indwidth <= wQUAD;
  parwidth <= pBYTE;
  admode <= sPREINDIRECT;
when "0000000100" =>          -- $04, TSB Zeropage: zp  (cmos)
  operation <= xTSB;
  parwidth <= pw_bl;
  admode <= sABSOLUTE;
when "0000000101" =>          -- $05, ORA Zeropage: zp 
  operation <= xORA;
  parwidth <= pw_bl;
  admode <= sABSOLUTE;
when "0000000110" =>          -- $06, ASL Zeropage: zp 
  operation <= xASL;
  parwidth <= pw_bl;
  admode <= sABSOLUTE;
when "0000000111" =>          -- $07, JMP Absolute indirect 64bit: [[abs]]  (65k)
  operation <= xJMP;
  default_le <= eSIGN;
  indwidth <= wQUAD;
  parwidth <= pWORD;
  admode <= sINDIRECT;
when "0000001000" =>          -- $08, PHP Implied:  
  operation <= xPHP;
  admode <= sIMPLIED;
when "0000001001" =>          -- $09, ORA Immediate: #byte 
  operation <= xORA;
  parwidth <= pw_rs;
  admode <= sIMMEDIATE;
when "0000001010" =>          -- $0a, ASL Accumulator:  
  operation <= xASL_A;
  admode <= sIMPLIED;
when "0000001100" =>          -- $0c, TSB Absolute 16bit: abs  (cmos)
  operation <= xTSB;
  parwidth <= pw_wq;
  admode <= sABSOLUTE;
when "0000001101" =>          -- $0d, ORA Absolute 16bit: abs 
  operation <= xORA;
  parwidth <= pw_wq;
  admode <= sABSOLUTE;
when "0000001110" =>          -- $0e, ASL Absolute 16bit: abs 
  operation <= xASL;
  parwidth <= pw_wq;
  admode <= sABSOLUTE;
when "0000010000" =>          -- $10, BPL Relative: rel 
  operation <= xBPL;
  parwidth <= pw_rs;
  admode <= sREL;
when "0000010001" =>          -- $11, ORA Zeropage indirect 16bit indexed with Y: (zp),Y 
  operation <= xORA;
  idxreg <= iYR;
  indwidth <= wWORD;
  parwidth <= pBYTE;
  admode <= sPOSTINDIRECT;
when "0000010010" =>          -- $12, ORA Zeropage indirect 16bit: (zp)  (cmos)
  operation <= xORA;
  indwidth <= wWORD;
  parwidth <= pBYTE;
  admode <= sINDIRECT;
when "0000010011" =>          -- $13, ORA Zeropage indirect 64bit indexed with Y: [[zp]],Y  (65k)
  operation <= xORA;
  idxreg <= iYR;
  indwidth <= wQUAD;
  parwidth <= pBYTE;
  admode <= sPOSTINDIRECT;
when "0000010100" =>          -- $14, TRB Zeropage: zp  (cmos)
  operation <= xTRB;
  parwidth <= pw_bl;
  admode <= sABSOLUTE;
when "0000010101" =>          -- $15, ORA Zeropage indexed with X: zp,X 
  operation <= xORA;
  idxreg <= iXR;
  parwidth <= pw_bl;
  admode <= sABSOLUTEIND;
when "0000010110" =>          -- $16, ASL Zeropage indexed with X: zp,X 
  operation <= xASL;
  idxreg <= iXR;
  parwidth <= pw_bl;
  admode <= sABSOLUTEIND;
when "0000010111" =>          -- $17, ORA Zeropage indirect 64bit: [[zp]]  (65k)
  operation <= xORA;
  indwidth <= wQUAD;
  parwidth <= pBYTE;
  admode <= sINDIRECT;
when "0000011000" =>          -- $18, CLC Implied:  
  operation <= xCLC;
  admode <= sIMPLIED;
when "0000011001" =>          -- $19, ORA Absolute 16bit indexed with Y: abs,Y 
  operation <= xORA;
  idxreg <= iYR;
  parwidth <= pw_wq;
  admode <= sABSOLUTEIND;
when "0000011010" =>          -- $1a, INC Accumulator:   (cmos)
  operation <= xINC_A;
  admode <= sIMPLIED;
when "0000011100" =>          -- $1c, TRB Absolute 16bit: abs  (cmos)
  operation <= xTRB;
  parwidth <= pw_wq;
  admode <= sABSOLUTE;
when "0000011101" =>          -- $1d, ORA Absolute 16bit indexed with X: abs,X 
  operation <= xORA;
  idxreg <= iXR;
  parwidth <= pw_wq;
  admode <= sABSOLUTEIND;
when "0000011110" =>          -- $1e, ASL Absolute 16bit indexed with X: abs,X 
  operation <= xASL;
  idxreg <= iXR;
  parwidth <= pw_wq;
  admode <= sABSOLUTEIND;
when "0000011111" =>          -- $1f, ASL Absolute 16bit indexed with Y: abs,Y  (65k)
  operation <= xASL;
  idxreg <= iYR;
  parwidth <= pw_wq;
  admode <= sABSOLUTEIND;
when "0000100000" =>          -- $20, JSR Address: abs 
  operation <= xJSR;
  default_le <= eSIGN;
  parwidth <= pw_wq;
  admode <= sADDR;
when "0000100001" =>          -- $21, AND Zeropage indexed with X indirect 16bit: (zp,X) 
  operation <= xAND;
  idxreg <= iXR;
  indwidth <= wWORD;
  parwidth <= pBYTE;
  admode <= sPREINDIRECT;
when "0000100010" =>          -- $22, STA Zeropage indexed with Y: zp,Y  (65k)
  operation <= xSTA;
  idxreg <= iYR;
  parwidth <= pw_bl;
  admode <= sABSOLUTEIND;
when "0000100011" =>          -- $23, AND Zeropage indexed with X indirect 64bit: [[zp,X]]  (65k)
  operation <= xAND;
  idxreg <= iXR;
  indwidth <= wQUAD;
  parwidth <= pBYTE;
  admode <= sPREINDIRECT;
when "0000100100" =>          -- $24, BIT Zeropage: zp 
  operation <= xBIT;
  parwidth <= pw_bl;
  admode <= sABSOLUTE;
when "0000100101" =>          -- $25, AND Zeropage: zp 
  operation <= xAND;
  parwidth <= pw_bl;
  admode <= sABSOLUTE;
when "0000100110" =>          -- $26, ROL Zeropage: zp 
  operation <= xROL;
  parwidth <= pw_bl;
  admode <= sABSOLUTE;
when "0000100111" =>          -- $27, JMP Absolute indexed with X indirect 64bit: [[abs,X]]  (65k)
  operation <= xJMP;
  default_le <= eSIGN;
  idxreg <= iXR;
  indwidth <= wQUAD;
  parwidth <= pWORD;
  admode <= sPREINDIRECT;
when "0000101000" =>          -- $28, PLP Implied:  
  operation <= xPLP;
  admode <= sIMPLIED;
when "0000101001" =>          -- $29, AND Immediate: #byte 
  operation <= xAND;
  parwidth <= pw_rs;
  admode <= sIMMEDIATE;
when "0000101010" =>          -- $2a, ROL Accumulator:  
  operation <= xROL_A;
  admode <= sIMPLIED;
when "0000101100" =>          -- $2c, BIT Absolute 16bit: abs 
  operation <= xBIT;
  parwidth <= pw_wq;
  admode <= sABSOLUTE;
when "0000101101" =>          -- $2d, AND Absolute 16bit: abs 
  operation <= xAND;
  parwidth <= pw_wq;
  admode <= sABSOLUTE;
when "0000101110" =>          -- $2e, ROL Absolute 16bit: abs 
  operation <= xROL;
  parwidth <= pw_wq;
  admode <= sABSOLUTE;
when "0000110000" =>          -- $30, BMI Relative: rel 
  operation <= xBMI;
  parwidth <= pw_rs;
  admode <= sREL;
when "0000110001" =>          -- $31, AND Zeropage indirect 16bit indexed with Y: (zp),Y 
  operation <= xAND;
  idxreg <= iYR;
  indwidth <= wWORD;
  parwidth <= pBYTE;
  admode <= sPOSTINDIRECT;
when "0000110010" =>          -- $32, AND Zeropage indirect 16bit: (zp)  (cmos)
  operation <= xAND;
  indwidth <= wWORD;
  parwidth <= pBYTE;
  admode <= sINDIRECT;
when "0000110011" =>          -- $33, AND Zeropage indirect 64bit indexed with Y: [[zp]],Y  (65k)
  operation <= xAND;
  idxreg <= iYR;
  indwidth <= wQUAD;
  parwidth <= pBYTE;
  admode <= sPOSTINDIRECT;
when "0000110100" =>          -- $34, BIT Zeropage indexed with X: zp,X  (cmos)
  operation <= xBIT;
  idxreg <= iXR;
  parwidth <= pw_bl;
  admode <= sABSOLUTEIND;
when "0000110101" =>          -- $35, AND Zeropage indexed with X: zp,X 
  operation <= xAND;
  idxreg <= iXR;
  parwidth <= pw_bl;
  admode <= sABSOLUTEIND;
when "0000110110" =>          -- $36, ROL Zeropage indexed with X: zp,X 
  operation <= xROL;
  idxreg <= iXR;
  parwidth <= pw_bl;
  admode <= sABSOLUTEIND;
when "0000110111" =>          -- $37, AND Zeropage indirect 64bit: [[zp]]  (65k)
  operation <= xAND;
  indwidth <= wQUAD;
  parwidth <= pBYTE;
  admode <= sINDIRECT;
when "0000111000" =>          -- $38, SEC Implied:  
  operation <= xSEC;
  admode <= sIMPLIED;
when "0000111001" =>          -- $39, AND Absolute 16bit indexed with Y: abs,Y 
  operation <= xAND;
  idxreg <= iYR;
  parwidth <= pw_wq;
  admode <= sABSOLUTEIND;
when "0000111010" =>          -- $3a, DEC Accumulator:   (cmos)
  operation <= xDEC_A;
  admode <= sIMPLIED;
when "0000111100" =>          -- $3c, BIT Absolute 16bit indexed with X: abs,X  (cmos)
  operation <= xBIT;
  idxreg <= iXR;
  parwidth <= pw_wq;
  admode <= sABSOLUTEIND;
when "0000111101" =>          -- $3d, AND Absolute 16bit indexed with X: abs,X 
  operation <= xAND;
  idxreg <= iXR;
  parwidth <= pw_wq;
  admode <= sABSOLUTEIND;
when "0000111110" =>          -- $3e, ROL Absolute 16bit indexed with X: abs,X 
  operation <= xROL;
  idxreg <= iXR;
  parwidth <= pw_wq;
  admode <= sABSOLUTEIND;
when "0000111111" =>          -- $3f, ROL Absolute 16bit indexed with Y: abs,Y  (65k)
  operation <= xROL;
  idxreg <= iYR;
  parwidth <= pw_wq;
  admode <= sABSOLUTEIND;
when "0001000000" =>          -- $40, RTI Implied:  
  operation <= xRTI;
  admode <= sIMPLIED;
when "0001000001" =>          -- $41, EOR Zeropage indexed with X indirect 16bit: (zp,X) 
  operation <= xEOR;
  idxreg <= iXR;
  indwidth <= wWORD;
  parwidth <= pBYTE;
  admode <= sPREINDIRECT;
when "0001000010" =>          -- $42, LDA Absolute indirect 16bit indexed with Y: (abs),Y  (65k)
  operation <= xLDA;
  default_le <= eZERO;
  idxreg <= iYR;
  indwidth <= wWORD;
  parwidth <= pWORD;
  admode <= sPOSTINDIRECT;
when "0001000011" =>          -- $43, EOR Zeropage indexed with X indirect 64bit: [[zp,X]]  (65k)
  operation <= xEOR;
  idxreg <= iXR;
  indwidth <= wQUAD;
  parwidth <= pBYTE;
  admode <= sPREINDIRECT;
when "0001000100" =>          -- $44, BSR Relative 16bit (BSR): relwide  (65k)
  operation <= xBSR;
  parwidth <= pw_wq;
  admode <= sREL;
when "0001000101" =>          -- $45, EOR Zeropage: zp 
  operation <= xEOR;
  parwidth <= pw_bl;
  admode <= sABSOLUTE;
when "0001000110" =>          -- $46, LSR Zeropage: zp 
  operation <= xLSR;
  parwidth <= pw_bl;
  admode <= sABSOLUTE;
when "0001000111" =>          -- $47, LDA Absolute indirect 64bit indexed with Y: [[abs]],Y  (65k)
  operation <= xLDA;
  default_le <= eZERO;
  idxreg <= iYR;
  indwidth <= wQUAD;
  parwidth <= pWORD;
  admode <= sPOSTINDIRECT;
when "0001001000" =>          -- $48, PHA Implied:  
  operation <= xPHA;
  admode <= sIMPLIED;
when "0001001001" =>          -- $49, EOR Immediate: #byte 
  operation <= xEOR;
  parwidth <= pw_rs;
  admode <= sIMMEDIATE;
when "0001001010" =>          -- $4a, LSR Accumulator:  
  operation <= xLSR_A;
  admode <= sIMPLIED;
when "0001001100" =>          -- $4c, JMP Address: abs 
  operation <= xJMP;
  default_le <= eSIGN;
  parwidth <= pw_wq;
  admode <= sADDR;
when "0001001101" =>          -- $4d, EOR Absolute 16bit: abs 
  operation <= xEOR;
  parwidth <= pw_wq;
  admode <= sABSOLUTE;
when "0001001110" =>          -- $4e, LSR Absolute 16bit: abs 
  operation <= xLSR;
  parwidth <= pw_wq;
  admode <= sABSOLUTE;
when "0001010000" =>          -- $50, BVC Relative: rel 
  operation <= xBVC;
  parwidth <= pw_rs;
  admode <= sREL;
when "0001010001" =>          -- $51, EOR Zeropage indirect 16bit indexed with Y: (zp),Y 
  operation <= xEOR;
  idxreg <= iYR;
  indwidth <= wWORD;
  parwidth <= pBYTE;
  admode <= sPOSTINDIRECT;
when "0001010010" =>          -- $52, EOR Zeropage indirect 16bit: (zp)  (cmos)
  operation <= xEOR;
  indwidth <= wWORD;
  parwidth <= pBYTE;
  admode <= sINDIRECT;
when "0001010011" =>          -- $53, EOR Zeropage indirect 64bit indexed with Y: [[zp]],Y  (65k)
  operation <= xEOR;
  idxreg <= iYR;
  indwidth <= wQUAD;
  parwidth <= pBYTE;
  admode <= sPOSTINDIRECT;
when "0001010101" =>          -- $55, EOR Zeropage indexed with X: zp,X 
  operation <= xEOR;
  idxreg <= iXR;
  parwidth <= pw_bl;
  admode <= sABSOLUTEIND;
when "0001010110" =>          -- $56, LSR Zeropage indexed with X: zp,X 
  operation <= xLSR;
  idxreg <= iXR;
  parwidth <= pw_bl;
  admode <= sABSOLUTEIND;
when "0001010111" =>          -- $57, EOR Zeropage indirect 64bit: [[zp]]  (65k)
  operation <= xEOR;
  indwidth <= wQUAD;
  parwidth <= pBYTE;
  admode <= sINDIRECT;
when "0001011000" =>          -- $58, CLI Implied:  
  operation <= xCLI;
  admode <= sIMPLIED;
when "0001011001" =>          -- $59, EOR Absolute 16bit indexed with Y: abs,Y 
  operation <= xEOR;
  idxreg <= iYR;
  parwidth <= pw_wq;
  admode <= sABSOLUTEIND;
when "0001011010" =>          -- $5a, PHY Implied:   (cmos)
  operation <= xPHY;
  admode <= sIMPLIED;
when "0001011101" =>          -- $5d, EOR Absolute 16bit indexed with X: abs,X 
  operation <= xEOR;
  idxreg <= iXR;
  parwidth <= pw_wq;
  admode <= sABSOLUTEIND;
when "0001011110" =>          -- $5e, LSR Absolute 16bit indexed with X: abs,X 
  operation <= xLSR;
  idxreg <= iXR;
  parwidth <= pw_wq;
  admode <= sABSOLUTEIND;
when "0001011111" =>          -- $5f, LSR Absolute 16bit indexed with Y: abs,Y  (65k)
  operation <= xLSR;
  idxreg <= iYR;
  parwidth <= pw_wq;
  admode <= sABSOLUTEIND;
when "0001100000" =>          -- $60, RTS Implied:  
  operation <= xRTS;
  admode <= sIMPLIED;
when "0001100001" =>          -- $61, ADC Zeropage indexed with X indirect 16bit: (zp,X) 
  operation <= xADC;
  idxreg <= iXR;
  indwidth <= wWORD;
  parwidth <= pBYTE;
  admode <= sPREINDIRECT;
when "0001100010" =>          -- $62, LDA Absolute indexed with X indirect 16bit: (abs,X)  (65k)
  operation <= xLDA;
  default_le <= eZERO;
  idxreg <= iXR;
  indwidth <= wWORD;
  parwidth <= pWORD;
  admode <= sPREINDIRECT;
when "0001100011" =>          -- $63, ADC Zeropage indexed with X indirect 64bit: [[zp,X]]  (65k)
  operation <= xADC;
  idxreg <= iXR;
  indwidth <= wQUAD;
  parwidth <= pBYTE;
  admode <= sPREINDIRECT;
when "0001100100" =>          -- $64, STZ Zeropage: zp  (cmos)
  operation <= xSTZ;
  parwidth <= pw_bl;
  admode <= sABSOLUTE;
when "0001100101" =>          -- $65, ADC Zeropage: zp 
  operation <= xADC;
  parwidth <= pw_bl;
  admode <= sABSOLUTE;
when "0001100110" =>          -- $66, ROR Zeropage: zp 
  operation <= xROR;
  parwidth <= pw_bl;
  admode <= sABSOLUTE;
when "0001100111" =>          -- $67, LDA Absolute indexed with X indirect 64bit: [[abs,X]]  (65k)
  operation <= xLDA;
  default_le <= eZERO;
  idxreg <= iXR;
  indwidth <= wQUAD;
  parwidth <= pWORD;
  admode <= sPREINDIRECT;
when "0001101000" =>          -- $68, PLA Implied:  
  operation <= xPLA;
  admode <= sIMPLIED;
when "0001101001" =>          -- $69, ADC Immediate: #byte 
  operation <= xADC;
  parwidth <= pw_rs;
  admode <= sIMMEDIATE;
when "0001101010" =>          -- $6a, ROR Accumulator:  
  operation <= xROR_A;
  admode <= sIMPLIED;
when "0001101100" =>          -- $6c, JMP Absolute indirect 16bit: (abs) 
  operation <= xJMP;
  default_le <= eSIGN;
  indwidth <= wWORD;
  parwidth <= pWORD;
  admode <= sINDIRECT;
when "0001101101" =>          -- $6d, ADC Absolute 16bit: abs 
  operation <= xADC;
  parwidth <= pw_wq;
  admode <= sABSOLUTE;
when "0001101110" =>          -- $6e, ROR Absolute 16bit: abs 
  operation <= xROR;
  parwidth <= pw_wq;
  admode <= sABSOLUTE;
when "0001110000" =>          -- $70, BVS Relative: rel 
  operation <= xBVS;
  parwidth <= pw_rs;
  admode <= sREL;
when "0001110001" =>          -- $71, ADC Zeropage indirect 16bit indexed with Y: (zp),Y 
  operation <= xADC;
  idxreg <= iYR;
  indwidth <= wWORD;
  parwidth <= pBYTE;
  admode <= sPOSTINDIRECT;
when "0001110010" =>          -- $72, ADC Zeropage indirect 16bit: (zp)  (cmos)
  operation <= xADC;
  indwidth <= wWORD;
  parwidth <= pBYTE;
  admode <= sINDIRECT;
when "0001110011" =>          -- $73, ADC Zeropage indirect 64bit indexed with Y: [[zp]],Y  (65k)
  operation <= xADC;
  idxreg <= iYR;
  indwidth <= wQUAD;
  parwidth <= pBYTE;
  admode <= sPOSTINDIRECT;
when "0001110100" =>          -- $74, STZ Zeropage indexed with X: zp,X  (cmos)
  operation <= xSTZ;
  idxreg <= iXR;
  parwidth <= pw_bl;
  admode <= sABSOLUTEIND;
when "0001110101" =>          -- $75, ADC Zeropage indexed with X: zp,X 
  operation <= xADC;
  idxreg <= iXR;
  parwidth <= pw_bl;
  admode <= sABSOLUTEIND;
when "0001110110" =>          -- $76, ROR Zeropage indexed with X: zp,X 
  operation <= xROR;
  idxreg <= iXR;
  parwidth <= pw_bl;
  admode <= sABSOLUTEIND;
when "0001110111" =>          -- $77, ADC Zeropage indirect 64bit: [[zp]]  (65k)
  operation <= xADC;
  indwidth <= wQUAD;
  parwidth <= pBYTE;
  admode <= sINDIRECT;
when "0001111000" =>          -- $78, SEI Implied:  
  operation <= xSEI;
  admode <= sIMPLIED;
when "0001111001" =>          -- $79, ADC Absolute 16bit indexed with Y: abs,Y 
  operation <= xADC;
  idxreg <= iYR;
  parwidth <= pw_wq;
  admode <= sABSOLUTEIND;
when "0001111010" =>          -- $7a, PLY Implied:   (cmos)
  operation <= xPLY;
  admode <= sIMPLIED;
when "0001111100" =>          -- $7c, JMP Absolute indexed with X indirect 16bit: (abs,X)  (cmos)
  operation <= xJMP;
  default_le <= eSIGN;
  idxreg <= iXR;
  indwidth <= wWORD;
  parwidth <= pWORD;
  admode <= sPREINDIRECT;
when "0001111101" =>          -- $7d, ADC Absolute 16bit indexed with X: abs,X 
  operation <= xADC;
  idxreg <= iXR;
  parwidth <= pw_wq;
  admode <= sABSOLUTEIND;
when "0001111110" =>          -- $7e, ROR Absolute 16bit indexed with X: abs,X 
  operation <= xROR;
  idxreg <= iXR;
  parwidth <= pw_wq;
  admode <= sABSOLUTEIND;
when "0001111111" =>          -- $7f, ROR Absolute 16bit indexed with Y: abs,Y  (65k)
  operation <= xROR;
  idxreg <= iYR;
  parwidth <= pw_wq;
  admode <= sABSOLUTEIND;
when "0010000000" =>          -- $80, BRA Relative: rel  (cmos)
  operation <= xBRA;
  parwidth <= pw_rs;
  admode <= sREL;
when "0010000001" =>          -- $81, STA Zeropage indexed with X indirect 16bit: (zp,X) 
  operation <= xSTA;
  idxreg <= iXR;
  indwidth <= wWORD;
  parwidth <= pBYTE;
  admode <= sPREINDIRECT;
when "0010000010" =>          -- $82, BSR Relative (BSR): rel  (65k)
  operation <= xBSR;
  parwidth <= pw_bl;
  admode <= sREL;
when "0010000011" =>          -- $83, STA Zeropage indexed with X indirect 64bit: [[zp,X]]  (65k)
  operation <= xSTA;
  idxreg <= iXR;
  indwidth <= wQUAD;
  parwidth <= pBYTE;
  admode <= sPREINDIRECT;
when "0010000100" =>          -- $84, STY Zeropage: zp 
  operation <= xSTY;
  parwidth <= pw_bl;
  admode <= sABSOLUTE;
when "0010000101" =>          -- $85, STA Zeropage: zp 
  operation <= xSTA;
  parwidth <= pw_bl;
  admode <= sABSOLUTE;
when "0010000110" =>          -- $86, STX Zeropage: zp 
  operation <= xSTX;
  parwidth <= pw_bl;
  admode <= sABSOLUTE;
when "0010000111" =>          -- $87, JSR Absolute indirect 64bit: [[abs]]  (65k)
  operation <= xJSR;
  default_le <= eSIGN;
  indwidth <= wQUAD;
  parwidth <= pWORD;
  admode <= sINDIRECT;
when "0010001000" =>          -- $88, DEY Implied:  
  operation <= xDEY;
  admode <= sIMPLIED;
when "0010001001" =>          -- $89, BIT Immediate: #byte  (cmos)
  operation <= xBIT;
  parwidth <= pw_rs;
  admode <= sIMMEDIATE;
when "0010001010" =>          -- $8a, TXA Implied:  
  operation <= xTXA;
  admode <= sIMPLIED;
when "0010001100" =>          -- $8c, STY Absolute 16bit: abs 
  operation <= xSTY;
  parwidth <= pw_wq;
  admode <= sABSOLUTE;
when "0010001101" =>          -- $8d, STA Absolute 16bit: abs 
  operation <= xSTA;
  parwidth <= pw_wq;
  admode <= sABSOLUTE;
when "0010001110" =>          -- $8e, STX Absolute 16bit: abs 
  operation <= xSTX;
  parwidth <= pw_wq;
  admode <= sABSOLUTE;
when "0010010000" =>          -- $90, BCC Relative: rel 
  operation <= xBCC;
  parwidth <= pw_rs;
  admode <= sREL;
when "0010010001" =>          -- $91, STA Zeropage indirect 16bit indexed with Y: (zp),Y 
  operation <= xSTA;
  idxreg <= iYR;
  indwidth <= wWORD;
  parwidth <= pBYTE;
  admode <= sPOSTINDIRECT;
when "0010010010" =>          -- $92, STA Zeropage indirect 16bit: (zp)  (cmos)
  operation <= xSTA;
  indwidth <= wWORD;
  parwidth <= pBYTE;
  admode <= sINDIRECT;
when "0010010011" =>          -- $93, STA Zeropage indirect 64bit indexed with Y: [[zp]],Y  (65k)
  operation <= xSTA;
  idxreg <= iYR;
  indwidth <= wQUAD;
  parwidth <= pBYTE;
  admode <= sPOSTINDIRECT;
when "0010010100" =>          -- $94, STY Zeropage indexed with X: zp,X 
  operation <= xSTY;
  idxreg <= iXR;
  parwidth <= pw_bl;
  admode <= sABSOLUTEIND;
when "0010010101" =>          -- $95, STA Zeropage indexed with X: zp,X 
  operation <= xSTA;
  idxreg <= iXR;
  parwidth <= pw_bl;
  admode <= sABSOLUTEIND;
when "0010010110" =>          -- $96, STX Zeropage indexed with Y: zp,Y 
  operation <= xSTX;
  idxreg <= iYR;
  parwidth <= pw_bl;
  admode <= sABSOLUTEIND;
when "0010010111" =>          -- $97, STA Zeropage indirect 64bit: [[zp]]  (65k)
  operation <= xSTA;
  indwidth <= wQUAD;
  parwidth <= pBYTE;
  admode <= sINDIRECT;
when "0010011000" =>          -- $98, TYA Implied:  
  operation <= xTYA;
  admode <= sIMPLIED;
when "0010011001" =>          -- $99, STA Absolute 16bit indexed with Y: abs,Y 
  operation <= xSTA;
  idxreg <= iYR;
  parwidth <= pw_wq;
  admode <= sABSOLUTEIND;
when "0010011010" =>          -- $9a, TXS Implied:  
  operation <= xTXS;
  admode <= sIMPLIED;
when "0010011100" =>          -- $9c, STZ Absolute 16bit: abs  (cmos)
  operation <= xSTZ;
  parwidth <= pw_wq;
  admode <= sABSOLUTE;
when "0010011101" =>          -- $9d, STA Absolute 16bit indexed with X: abs,X 
  operation <= xSTA;
  idxreg <= iXR;
  parwidth <= pw_wq;
  admode <= sABSOLUTEIND;
when "0010011110" =>          -- $9e, STZ Absolute 16bit indexed with X: abs,X  (cmos)
  operation <= xSTZ;
  idxreg <= iXR;
  parwidth <= pw_wq;
  admode <= sABSOLUTEIND;
when "0010011111" =>          -- $9f, STY Absolute 16bit indexed with X: abs,X  (65k)
  operation <= xSTY;
  idxreg <= iXR;
  parwidth <= pw_wq;
  admode <= sABSOLUTEIND;
when "0010100000" =>          -- $a0, LDY Immediate: #byte 
  operation <= xLDY;
  default_le <= eZERO;
  parwidth <= pw_rs;
  admode <= sIMMEDIATE;
when "0010100001" =>          -- $a1, LDA Zeropage indexed with X indirect 16bit: (zp,X) 
  operation <= xLDA;
  default_le <= eZERO;
  idxreg <= iXR;
  indwidth <= wWORD;
  parwidth <= pBYTE;
  admode <= sPREINDIRECT;
when "0010100010" =>          -- $a2, LDX Immediate: #byte 
  operation <= xLDX;
  default_le <= eZERO;
  parwidth <= pw_rs;
  admode <= sIMMEDIATE;
when "0010100011" =>          -- $a3, LDA Zeropage indexed with X indirect 64bit: [[zp,X]]  (65k)
  operation <= xLDA;
  default_le <= eZERO;
  idxreg <= iXR;
  indwidth <= wQUAD;
  parwidth <= pBYTE;
  admode <= sPREINDIRECT;
when "0010100100" =>          -- $a4, LDY Zeropage: zp 
  operation <= xLDY;
  default_le <= eZERO;
  parwidth <= pw_bl;
  admode <= sABSOLUTE;
when "0010100101" =>          -- $a5, LDA Zeropage: zp 
  operation <= xLDA;
  default_le <= eZERO;
  parwidth <= pw_bl;
  admode <= sABSOLUTE;
when "0010100110" =>          -- $a6, LDX Zeropage: zp 
  operation <= xLDX;
  default_le <= eZERO;
  parwidth <= pw_bl;
  admode <= sABSOLUTE;
when "0010100111" =>          -- $a7, JSR Absolute indexed with X indirect 64bit: [[abs,X]]  (65k)
  operation <= xJSR;
  default_le <= eSIGN;
  idxreg <= iXR;
  indwidth <= wQUAD;
  parwidth <= pWORD;
  admode <= sPREINDIRECT;
when "0010101000" =>          -- $a8, TAY Implied:  
  operation <= xTAY;
  admode <= sIMPLIED;
when "0010101001" =>          -- $a9, LDA Immediate: #byte 
  operation <= xLDA;
  default_le <= eZERO;
  parwidth <= pw_rs;
  admode <= sIMMEDIATE;
when "0010101010" =>          -- $aa, TAX Implied:  
  operation <= xTAX;
  admode <= sIMPLIED;
when "0010101100" =>          -- $ac, LDY Absolute 16bit: abs 
  operation <= xLDY;
  default_le <= eZERO;
  parwidth <= pw_wq;
  admode <= sABSOLUTE;
when "0010101101" =>          -- $ad, LDA Absolute 16bit: abs 
  operation <= xLDA;
  default_le <= eZERO;
  parwidth <= pw_wq;
  admode <= sABSOLUTE;
when "0010101110" =>          -- $ae, LDX Absolute 16bit: abs 
  operation <= xLDX;
  default_le <= eZERO;
  parwidth <= pw_wq;
  admode <= sABSOLUTE;
when "0010110000" =>          -- $b0, BCS Relative: rel 
  operation <= xBCS;
  parwidth <= pw_rs;
  admode <= sREL;
when "0010110001" =>          -- $b1, LDA Zeropage indirect 16bit indexed with Y: (zp),Y 
  operation <= xLDA;
  default_le <= eZERO;
  idxreg <= iYR;
  indwidth <= wWORD;
  parwidth <= pBYTE;
  admode <= sPOSTINDIRECT;
when "0010110010" =>          -- $b2, LDA Zeropage indirect 16bit: (zp)  (cmos)
  operation <= xLDA;
  default_le <= eZERO;
  indwidth <= wWORD;
  parwidth <= pBYTE;
  admode <= sINDIRECT;
when "0010110011" =>          -- $b3, LDA Zeropage indirect 64bit indexed with Y: [[zp]],Y  (65k)
  operation <= xLDA;
  default_le <= eZERO;
  idxreg <= iYR;
  indwidth <= wQUAD;
  parwidth <= pBYTE;
  admode <= sPOSTINDIRECT;
when "0010110100" =>          -- $b4, LDY Zeropage indexed with X: zp,X 
  operation <= xLDY;
  default_le <= eZERO;
  idxreg <= iXR;
  parwidth <= pw_bl;
  admode <= sABSOLUTEIND;
when "0010110101" =>          -- $b5, LDA Zeropage indexed with X: zp,X 
  operation <= xLDA;
  default_le <= eZERO;
  idxreg <= iXR;
  parwidth <= pw_bl;
  admode <= sABSOLUTEIND;
when "0010110110" =>          -- $b6, LDX Zeropage indexed with Y: zp,Y 
  operation <= xLDX;
  default_le <= eZERO;
  idxreg <= iYR;
  parwidth <= pw_bl;
  admode <= sABSOLUTEIND;
when "0010110111" =>          -- $b7, LDA Zeropage indirect 64bit: [[zp]]  (65k)
  operation <= xLDA;
  default_le <= eZERO;
  indwidth <= wQUAD;
  parwidth <= pBYTE;
  admode <= sINDIRECT;
when "0010111000" =>          -- $b8, CLV Implied:  
  operation <= xCLV;
  admode <= sIMPLIED;
when "0010111001" =>          -- $b9, LDA Absolute 16bit indexed with Y: abs,Y 
  operation <= xLDA;
  default_le <= eZERO;
  idxreg <= iYR;
  parwidth <= pw_wq;
  admode <= sABSOLUTEIND;
when "0010111010" =>          -- $ba, TSX Implied:  
  operation <= xTSX;
  admode <= sIMPLIED;
when "0010111100" =>          -- $bc, LDY Absolute 16bit indexed with X: abs,X 
  operation <= xLDY;
  default_le <= eZERO;
  idxreg <= iXR;
  parwidth <= pw_wq;
  admode <= sABSOLUTEIND;
when "0010111101" =>          -- $bd, LDA Absolute 16bit indexed with X: abs,X 
  operation <= xLDA;
  default_le <= eZERO;
  idxreg <= iXR;
  parwidth <= pw_wq;
  admode <= sABSOLUTEIND;
when "0010111110" =>          -- $be, LDX Absolute 16bit indexed with Y: abs,Y 
  operation <= xLDX;
  default_le <= eZERO;
  idxreg <= iYR;
  parwidth <= pw_wq;
  admode <= sABSOLUTEIND;
when "0010111111" =>          -- $bf, STX Absolute 16bit indexed with Y: abs,Y  (65k)
  operation <= xSTX;
  idxreg <= iYR;
  parwidth <= pw_wq;
  admode <= sABSOLUTEIND;
when "0011000000" =>          -- $c0, CPY Immediate: #byte 
  operation <= xCPY;
  parwidth <= pw_rs;
  admode <= sIMMEDIATE;
when "0011000001" =>          -- $c1, CMP Zeropage indexed with X indirect 16bit: (zp,X) 
  operation <= xCMP;
  idxreg <= iXR;
  indwidth <= wWORD;
  parwidth <= pBYTE;
  admode <= sPREINDIRECT;
when "0011000010" =>          -- $c2, STA Absolute indirect 16bit indexed with Y: (abs),Y  (65k)
  operation <= xSTA;
  idxreg <= iYR;
  indwidth <= wWORD;
  parwidth <= pWORD;
  admode <= sPOSTINDIRECT;
when "0011000011" =>          -- $c3, CMP Zeropage indexed with X indirect 64bit: [[zp,X]]  (65k)
  operation <= xCMP;
  idxreg <= iXR;
  indwidth <= wQUAD;
  parwidth <= pBYTE;
  admode <= sPREINDIRECT;
when "0011000100" =>          -- $c4, CPY Zeropage: zp 
  operation <= xCPY;
  parwidth <= pw_bl;
  admode <= sABSOLUTE;
when "0011000101" =>          -- $c5, CMP Zeropage: zp 
  operation <= xCMP;
  parwidth <= pw_bl;
  admode <= sABSOLUTE;
when "0011000110" =>          -- $c6, DEC Zeropage: zp 
  operation <= xDEC;
  parwidth <= pw_bl;
  admode <= sABSOLUTE;
when "0011000111" =>          -- $c7, STA Absolute indirect 64bit indexed with Y: [[abs]],Y  (65k)
  operation <= xSTA;
  idxreg <= iYR;
  indwidth <= wQUAD;
  parwidth <= pWORD;
  admode <= sPOSTINDIRECT;
when "0011001000" =>          -- $c8, INY Implied:  
  operation <= xINY;
  admode <= sIMPLIED;
when "0011001001" =>          -- $c9, CMP Immediate: #byte 
  operation <= xCMP;
  parwidth <= pw_rs;
  admode <= sIMMEDIATE;
when "0011001010" =>          -- $ca, DEX Implied:  
  operation <= xDEX;
  admode <= sIMPLIED;
when "0011001100" =>          -- $cc, CPY Absolute 16bit: abs 
  operation <= xCPY;
  parwidth <= pw_wq;
  admode <= sABSOLUTE;
when "0011001101" =>          -- $cd, CMP Absolute 16bit: abs 
  operation <= xCMP;
  parwidth <= pw_wq;
  admode <= sABSOLUTE;
when "0011001110" =>          -- $ce, DEC Absolute 16bit: abs 
  operation <= xDEC;
  parwidth <= pw_wq;
  admode <= sABSOLUTE;
when "0011010000" =>          -- $d0, BNE Relative: rel 
  operation <= xBNE;
  parwidth <= pw_rs;
  admode <= sREL;
when "0011010001" =>          -- $d1, CMP Zeropage indirect 16bit indexed with Y: (zp),Y 
  operation <= xCMP;
  idxreg <= iYR;
  indwidth <= wWORD;
  parwidth <= pBYTE;
  admode <= sPOSTINDIRECT;
when "0011010010" =>          -- $d2, CMP Zeropage indirect 16bit: (zp)  (cmos)
  operation <= xCMP;
  indwidth <= wWORD;
  parwidth <= pBYTE;
  admode <= sINDIRECT;
when "0011010011" =>          -- $d3, CMP Zeropage indirect 64bit indexed with Y: [[zp]],Y  (65k)
  operation <= xCMP;
  idxreg <= iYR;
  indwidth <= wQUAD;
  parwidth <= pBYTE;
  admode <= sPOSTINDIRECT;
when "0011010101" =>          -- $d5, CMP Zeropage indexed with X: zp,X 
  operation <= xCMP;
  idxreg <= iXR;
  parwidth <= pw_bl;
  admode <= sABSOLUTEIND;
when "0011010110" =>          -- $d6, DEC Zeropage indexed with X: zp,X 
  operation <= xDEC;
  idxreg <= iXR;
  parwidth <= pw_bl;
  admode <= sABSOLUTEIND;
when "0011010111" =>          -- $d7, CMP Zeropage indirect 64bit: [[zp]]  (65k)
  operation <= xCMP;
  indwidth <= wQUAD;
  parwidth <= pBYTE;
  admode <= sINDIRECT;
when "0011011000" =>          -- $d8, CLD Implied:  
  operation <= xCLD;
  admode <= sIMPLIED;
when "0011011001" =>          -- $d9, CMP Absolute 16bit indexed with Y: abs,Y 
  operation <= xCMP;
  idxreg <= iYR;
  parwidth <= pw_wq;
  admode <= sABSOLUTEIND;
when "0011011010" =>          -- $da, PHX Implied:   (cmos)
  operation <= xPHX;
  admode <= sIMPLIED;
when "0011011100" =>          -- $dc, JSR Absolute indirect 16bit: (abs)  (65k)
  operation <= xJSR;
  default_le <= eSIGN;
  indwidth <= wWORD;
  parwidth <= pWORD;
  admode <= sINDIRECT;
when "0011011101" =>          -- $dd, CMP Absolute 16bit indexed with X: abs,X 
  operation <= xCMP;
  idxreg <= iXR;
  parwidth <= pw_wq;
  admode <= sABSOLUTEIND;
when "0011011110" =>          -- $de, DEC Absolute 16bit indexed with X: abs,X 
  operation <= xDEC;
  idxreg <= iXR;
  parwidth <= pw_wq;
  admode <= sABSOLUTEIND;
when "0011011111" =>          -- $df, DEC Absolute 16bit indexed with Y: abs,Y  (65k)
  operation <= xDEC;
  idxreg <= iYR;
  parwidth <= pw_wq;
  admode <= sABSOLUTEIND;
when "0011100000" =>          -- $e0, CPX Immediate: #byte 
  operation <= xCPX;
  parwidth <= pw_rs;
  admode <= sIMMEDIATE;
when "0011100001" =>          -- $e1, SBC Zeropage indexed with X indirect 16bit: (zp,X) 
  operation <= xSBC;
  idxreg <= iXR;
  indwidth <= wWORD;
  parwidth <= pBYTE;
  admode <= sPREINDIRECT;
when "0011100010" =>          -- $e2, STA Absolute indexed with X indirect 16bit: (abs,X)  (65k)
  operation <= xSTA;
  idxreg <= iXR;
  indwidth <= wWORD;
  parwidth <= pWORD;
  admode <= sPREINDIRECT;
when "0011100011" =>          -- $e3, SBC Zeropage indexed with X indirect 64bit: [[zp,X]]  (65k)
  operation <= xSBC;
  idxreg <= iXR;
  indwidth <= wQUAD;
  parwidth <= pBYTE;
  admode <= sPREINDIRECT;
when "0011100100" =>          -- $e4, CPX Zeropage: zp 
  operation <= xCPX;
  parwidth <= pw_bl;
  admode <= sABSOLUTE;
when "0011100101" =>          -- $e5, SBC Zeropage: zp 
  operation <= xSBC;
  parwidth <= pw_bl;
  admode <= sABSOLUTE;
when "0011100110" =>          -- $e6, INC Zeropage: zp 
  operation <= xINC;
  parwidth <= pw_bl;
  admode <= sABSOLUTE;
when "0011100111" =>          -- $e7, STA Absolute indexed with X indirect 64bit: [[abs,X]]  (65k)
  operation <= xSTA;
  idxreg <= iXR;
  indwidth <= wQUAD;
  parwidth <= pWORD;
  admode <= sPREINDIRECT;
when "0011101000" =>          -- $e8, INX Implied:  
  operation <= xINX;
  admode <= sIMPLIED;
when "0011101001" =>          -- $e9, SBC Immediate: #byte 
  operation <= xSBC;
  parwidth <= pw_rs;
  admode <= sIMMEDIATE;
when "0011101010" =>          -- $ea, NOP Implied:  
  operation <= xNOP;
  admode <= sIMPLIED;
when "0011101100" =>          -- $ec, CPX Absolute 16bit: abs 
  operation <= xCPX;
  parwidth <= pw_wq;
  admode <= sABSOLUTE;
when "0011101101" =>          -- $ed, SBC Absolute 16bit: abs 
  operation <= xSBC;
  parwidth <= pw_wq;
  admode <= sABSOLUTE;
when "0011101110" =>          -- $ee, INC Absolute 16bit: abs 
  operation <= xINC;
  parwidth <= pw_wq;
  admode <= sABSOLUTE;
when "0011110000" =>          -- $f0, BEQ Relative: rel 
  operation <= xBEQ;
  parwidth <= pw_rs;
  admode <= sREL;
when "0011110001" =>          -- $f1, SBC Zeropage indirect 16bit indexed with Y: (zp),Y 
  operation <= xSBC;
  idxreg <= iYR;
  indwidth <= wWORD;
  parwidth <= pBYTE;
  admode <= sPOSTINDIRECT;
when "0011110010" =>          -- $f2, SBC Zeropage indirect 16bit: (zp)  (cmos)
  operation <= xSBC;
  indwidth <= wWORD;
  parwidth <= pBYTE;
  admode <= sINDIRECT;
when "0011110011" =>          -- $f3, SBC Zeropage indirect 64bit indexed with Y: [[zp]],Y  (65k)
  operation <= xSBC;
  idxreg <= iYR;
  indwidth <= wQUAD;
  parwidth <= pBYTE;
  admode <= sPOSTINDIRECT;
when "0011110100" =>          -- $f4, TRP Immediate: #byte  (65k)
  operation <= xTRP;
  parwidth <= pw_rs;
  admode <= sIMMEDIATE;
when "0011110101" =>          -- $f5, SBC Zeropage indexed with X: zp,X 
  operation <= xSBC;
  idxreg <= iXR;
  parwidth <= pw_bl;
  admode <= sABSOLUTEIND;
when "0011110110" =>          -- $f6, INC Zeropage indexed with X: zp,X 
  operation <= xINC;
  idxreg <= iXR;
  parwidth <= pw_bl;
  admode <= sABSOLUTEIND;
when "0011110111" =>          -- $f7, SBC Zeropage indirect 64bit: [[zp]]  (65k)
  operation <= xSBC;
  indwidth <= wQUAD;
  parwidth <= pBYTE;
  admode <= sINDIRECT;
when "0011111000" =>          -- $f8, SED Implied:  
  operation <= xSED;
  admode <= sIMPLIED;
when "0011111001" =>          -- $f9, SBC Absolute 16bit indexed with Y: abs,Y 
  operation <= xSBC;
  idxreg <= iYR;
  parwidth <= pw_wq;
  admode <= sABSOLUTEIND;
when "0011111010" =>          -- $fa, PLX Implied:   (cmos)
  operation <= xPLX;
  admode <= sIMPLIED;
when "0011111100" =>          -- $fc, JSR Absolute indexed with X indirect 16bit: (abs,X)  (65k)
  operation <= xJSR;
  default_le <= eSIGN;
  idxreg <= iXR;
  indwidth <= wWORD;
  parwidth <= pWORD;
  admode <= sPREINDIRECT;
when "0011111101" =>          -- $fd, SBC Absolute 16bit indexed with X: abs,X 
  operation <= xSBC;
  idxreg <= iXR;
  parwidth <= pw_wq;
  admode <= sABSOLUTEIND;
when "0011111110" =>          -- $fe, INC Absolute 16bit indexed with X: abs,X 
  operation <= xINC;
  idxreg <= iXR;
  parwidth <= pw_wq;
  admode <= sABSOLUTEIND;
when "0011111111" =>          -- $ff, INC Absolute 16bit indexed with Y: abs,Y  (65k)
  operation <= xINC;
  idxreg <= iYR;
  parwidth <= pw_wq;
  admode <= sABSOLUTEIND;
when "0100000010" =>          -- $02, LEA Zeropage indexed with Y: zp,Y  (65k)
  operation <= xLEA;
  idxreg <= iYR;
  parwidth <= pw_bl;
  admode <= sABSOLUTEIND;
when "0100000100" =>          -- $04, MVN Implied:   (65k)
  operation <= xMVN;
  admode <= sIMPLIED;
when "0100000110" =>          -- $06, ASR Zeropage: zp  (65k)
  operation <= xASR;
  parwidth <= pw_bl;
  admode <= sABSOLUTE;
when "0100001000" =>          -- $08, PHE Implied:   (65k)
  operation <= xPHE;
  admode <= sIMPLIED;
when "0100001001" =>          -- $09, ORA E indirect: (E)  (65k)
  operation <= xORA;
  admode <= sEINDIRECT;
when "0100001010" =>          -- $0a, ASR Accumulator:   (65k)
  operation <= xASR_A;
  admode <= sIMPLIED;
when "0100001100" =>          -- $0c, TSB E indirect: (E)  (65k)
  operation <= xTSB;
  admode <= sEINDIRECT;
when "0100001101" =>          -- $0d, ASL E indirect: (E)  (65k)
  operation <= xASL;
  admode <= sEINDIRECT;
when "0100001110" =>          -- $0e, ASR Absolute 16bit: abs  (65k)
  operation <= xASR;
  parwidth <= pw_wq;
  admode <= sABSOLUTE;
when "0100010100" =>          -- $14, MVP Implied:   (65k)
  operation <= xMVP;
  admode <= sIMPLIED;
when "0100010110" =>          -- $16, ASR Zeropage indexed with X: zp,X  (65k)
  operation <= xASR;
  idxreg <= iXR;
  parwidth <= pw_bl;
  admode <= sABSOLUTEIND;
when "0100011100" =>          -- $1c, TRB E indirect: (E)  (65k)
  operation <= xTRB;
  admode <= sEINDIRECT;
when "0100011101" =>          -- $1d, ASR E indirect: (E)  (65k)
  operation <= xASR;
  admode <= sEINDIRECT;
when "0100011110" =>          -- $1e, ASR Absolute 16bit indexed with X: abs,X  (65k)
  operation <= xASR;
  idxreg <= iXR;
  parwidth <= pw_wq;
  admode <= sABSOLUTEIND;
when "0100011111" =>          -- $1f, ASR Absolute 16bit indexed with Y: abs,Y  (65k)
  operation <= xASR;
  idxreg <= iYR;
  parwidth <= pw_wq;
  admode <= sABSOLUTEIND;
when "0100100000" =>          -- $20, JSR E indirect: (E)  (65k)
  operation <= xJSR;
  default_le <= eSIGN;
  admode <= sEINDIRECT;
when "0100100010" =>          -- $22, PEA Zeropage indexed with Y: zp,Y  (65k)
  operation <= xPEA;
  idxreg <= iYR;
  parwidth <= pw_bl;
  admode <= sABSOLUTEIND;
when "0100100100" =>          -- $24, FIL Implied:   (65k)
  operation <= xFIL;
  admode <= sIMPLIED;
when "0100100101" =>          -- $25, ADE Immediate: #byte  (65k)
  operation <= xADE;
  parwidth <= pw_rs;
  admode <= sIMMEDIATE;
when "0100100110" =>          -- $26, RDL Zeropage: zp  (65k)
  operation <= xRDL;
  parwidth <= pw_bl;
  admode <= sABSOLUTE;
when "0100101000" =>          -- $28, PLE Implied:   (65k)
  operation <= xPLE;
  admode <= sIMPLIED;
when "0100101001" =>          -- $29, AND E indirect: (E)  (65k)
  operation <= xAND;
  admode <= sEINDIRECT;
when "0100101010" =>          -- $2a, RDL Accumulator:   (65k)
  operation <= xRDL_A;
  admode <= sIMPLIED;
when "0100101101" =>          -- $2d, ROL E indirect: (E)  (65k)
  operation <= xROL;
  admode <= sEINDIRECT;
when "0100101110" =>          -- $2e, RDL Absolute 16bit: abs  (65k)
  operation <= xRDL;
  parwidth <= pw_wq;
  admode <= sABSOLUTE;
when "0100110100" =>          -- $34, BIT Accumulator:  
  operation <= xBIT_A;
  admode <= sIMPLIED;
when "0100110101" =>          -- $35, ADE Accumulator:   (65k)
  operation <= xADE_A;
  admode <= sIMPLIED;
when "0100110110" =>          -- $36, RDL Zeropage indexed with X: zp,X  (65k)
  operation <= xRDL;
  idxreg <= iXR;
  parwidth <= pw_bl;
  admode <= sABSOLUTEIND;
when "0100111001" =>          -- $39, LDE Immediate: #byte  (65k)
  operation <= xLDE;
  default_le <= eSIGN;
  parwidth <= pw_rs;
  admode <= sIMMEDIATE;
when "0100111101" =>          -- $3d, RDL E indirect: (E)  (65k)
  operation <= xRDL;
  admode <= sEINDIRECT;
when "0100111110" =>          -- $3e, RDL Absolute 16bit indexed with X: abs,X  (65k)
  operation <= xRDL;
  idxreg <= iXR;
  parwidth <= pw_wq;
  admode <= sABSOLUTEIND;
when "0100111111" =>          -- $3f, RDL Absolute 16bit indexed with Y: abs,Y  (65k)
  operation <= xRDL;
  idxreg <= iYR;
  parwidth <= pw_wq;
  admode <= sABSOLUTEIND;
when "0101000010" =>          -- $42, LEA Absolute indirect 16bit indexed with Y: (abs),Y  (65k)
  operation <= xLEA;
  idxreg <= iYR;
  indwidth <= wWORD;
  parwidth <= pWORD;
  admode <= sPOSTINDIRECT;
when "0101000100" =>          -- $44, LEA Relative 16bit: relwide  (65k)
  operation <= xLEA;
  parwidth <= pw_wq;
  admode <= sREL;
when "0101000101" =>          -- $45, ADS Immediate: #byte  (65k)
  operation <= xADS;
  parwidth <= pw_rs;
  admode <= sIMMEDIATE;
when "0101000110" =>          -- $46, LEA Zeropage: zp  (65k)
  operation <= xLEA;
  parwidth <= pw_bl;
  admode <= sABSOLUTE;
when "0101001000" =>          -- $48, PHB Implied:   (65k)
  operation <= xPHB;
  admode <= sIMPLIED;
when "0101001001" =>          -- $49, EOR E indirect: (E)  (65k)
  operation <= xEOR;
  admode <= sEINDIRECT;
when "0101001100" =>          -- $4c, JMP E indirect: (E)  (65k)
  operation <= xJMP;
  default_le <= eSIGN;
  admode <= sEINDIRECT;
when "0101001101" =>          -- $4d, LSR E indirect: (E)  (65k)
  operation <= xLSR;
  admode <= sEINDIRECT;
when "0101010100" =>          -- $54, PEA Relative 16bit: relwide  (65k)
  operation <= xPEA;
  parwidth <= pw_wq;
  admode <= sREL;
when "0101010101" =>          -- $55, ADS Accumulator:   (65k)
  operation <= xADS_A;
  admode <= sIMPLIED;
when "0101010110" =>          -- $56, LEA Zeropage indexed with X: zp,X  (65k)
  operation <= xLEA;
  idxreg <= iXR;
  parwidth <= pw_bl;
  admode <= sABSOLUTEIND;
when "0101011000" =>          -- $58, PRB Implied:   (65k)
  operation <= xPRB;
  admode <= sIMPLIED;
when "0101011001" =>          -- $59, LDB Immediate: #byte  (65k)
  operation <= xLDB;
  default_le <= eSIGN;
  parwidth <= pw_rs;
  admode <= sIMMEDIATE;
when "0101100010" =>          -- $62, LEA Absolute indexed with X indirect 16bit: (abs,X)  (65k)
  operation <= xLEA;
  idxreg <= iXR;
  indwidth <= wWORD;
  parwidth <= pWORD;
  admode <= sPREINDIRECT;
when "0101100100" =>          -- $64, RMB Implied:   (65k)
  operation <= xRMB;
  admode <= sIMPLIED;
when "0101100101" =>          -- $65, ADB Immediate: #byte  (65k)
  operation <= xADB;
  parwidth <= pw_rs;
  admode <= sIMMEDIATE;
when "0101100110" =>          -- $66, RDR Zeropage: zp 
  operation <= xRDR;
  parwidth <= pw_bl;
  admode <= sABSOLUTE;
when "0101101000" =>          -- $68, PLB Implied:   (65k)
  operation <= xPLB;
  admode <= sIMPLIED;
when "0101101001" =>          -- $69, ADC E indirect: (E)  (65k)
  operation <= xADC;
  admode <= sEINDIRECT;
when "0101101010" =>          -- $6a, RDR Accumulator:  
  operation <= xRDR_A;
  admode <= sIMPLIED;
when "0101101100" =>          -- $6c, JMP Address Long: long 
  operation <= xJMP;
  default_le <= eSIGN;
  parwidth <= pLONG;
  admode <= sADDR;
when "0101101101" =>          -- $6d, ROR E indirect: (E)  (65k)
  operation <= xROR;
  admode <= sEINDIRECT;
when "0101101110" =>          -- $6e, RDR Absolute 16bit: abs 
  operation <= xRDR;
  parwidth <= pw_wq;
  admode <= sABSOLUTE;
when "0101110100" =>          -- $74, WMB Implied:   (65k)
  operation <= xWMB;
  admode <= sIMPLIED;
when "0101110101" =>          -- $75, ADB Accumulator:   (65k)
  operation <= xADB_A;
  admode <= sIMPLIED;
when "0101110110" =>          -- $76, RDR Zeropage indexed with X: zp,X 
  operation <= xRDR;
  idxreg <= iXR;
  parwidth <= pw_bl;
  admode <= sABSOLUTEIND;
when "0101111101" =>          -- $7d, RDR E indirect: (E)  (65k)
  operation <= xRDR;
  admode <= sEINDIRECT;
when "0101111110" =>          -- $7e, RDR Absolute 16bit indexed with X: abs,X 
  operation <= xRDR;
  idxreg <= iXR;
  parwidth <= pw_wq;
  admode <= sABSOLUTEIND;
when "0101111111" =>          -- $7f, RDR Absolute 16bit indexed with Y: abs,Y 
  operation <= xRDR;
  idxreg <= iYR;
  parwidth <= pw_wq;
  admode <= sABSOLUTEIND;
when "0110000000" =>          -- $80, LEA Relative: rel  (65k)
  operation <= xLEA;
  parwidth <= pw_rs;
  admode <= sREL;
when "0110000001" =>          -- $81, PEA Zeropage indexed with X indirect 16bit: (zp,X)  (65k)
  operation <= xPEA;
  idxreg <= iXR;
  indwidth <= wWORD;
  parwidth <= pBYTE;
  admode <= sPREINDIRECT;
when "0110000010" =>          -- $82, PEA Relative: rel  (65k)
  operation <= xPEA;
  parwidth <= pw_rs;
  admode <= sREL;
when "0110000100" =>          -- $84, SCA E indirect: (E)  (65k)
  operation <= xSCA;
  admode <= sEINDIRECT;
when "0110000101" =>          -- $85, PEA Zeropage: zp  (65k)
  operation <= xPEA;
  parwidth <= pw_bl;
  admode <= sABSOLUTE;
when "0110001000" =>          -- $88, TAE Implied:   (65k)
  operation <= xTAE;
  admode <= sIMPLIED;
when "0110001001" =>          -- $89, BIT E indirect: (E)  (65k)
  operation <= xBIT;
  admode <= sEINDIRECT;
when "0110001010" =>          -- $8a, TYS Implied:   (65k)
  operation <= xTYS;
  admode <= sIMPLIED;
when "0110001100" =>          -- $8c, STY E indirect: (E)  (65k)
  operation <= xSTY;
  admode <= sEINDIRECT;
when "0110001101" =>          -- $8d, STA E indirect: (E)  (65k)
  operation <= xSTA;
  admode <= sEINDIRECT;
when "0110001110" =>          -- $8e, STX E indirect: (E)  (65k)
  operation <= xSTX;
  admode <= sEINDIRECT;
when "0110010001" =>          -- $91, PEA Zeropage indirect 16bit indexed with Y: (zp),Y  (65k)
  operation <= xPEA;
  idxreg <= iYR;
  indwidth <= wWORD;
  parwidth <= pBYTE;
  admode <= sPOSTINDIRECT;
when "0110010010" =>          -- $92, PEA Zeropage indirect 16bit: (zp)  (65k)
  operation <= xPEA;
  indwidth <= wWORD;
  parwidth <= pBYTE;
  admode <= sINDIRECT;
when "0110010100" =>          -- $94, LLA E indirect: (E)  (65k)
  operation <= xLLA;
  admode <= sEINDIRECT;
when "0110010101" =>          -- $95, PEA Zeropage indexed with X: zp,X  (65k)
  operation <= xPEA;
  idxreg <= iXR;
  parwidth <= pw_bl;
  admode <= sABSOLUTEIND;
when "0110011000" =>          -- $98, TEA Implied:   (65k)
  operation <= xTEA;
  admode <= sIMPLIED;
when "0110011001" =>          -- $99, PEA Absolute 16bit indexed with Y: abs,Y  (65k)
  operation <= xPEA;
  idxreg <= iYR;
  parwidth <= pw_wq;
  admode <= sABSOLUTEIND;
when "0110011010" =>          -- $9a, SXY Implied:   (65k)
  operation <= xSXY;
  admode <= sIMPLIED;
when "0110011100" =>          -- $9c, STZ E indirect: (E)  (65k)
  operation <= xSTZ;
  admode <= sEINDIRECT;
when "0110011110" =>          -- $9e, STZ Absolute 16bit indexed with Y: abs,Y  (65k)
  operation <= xSTZ;
  idxreg <= iYR;
  parwidth <= pw_wq;
  admode <= sABSOLUTEIND;
when "0110100000" =>          -- $a0, LDY E indirect: (E)  (65k)
  operation <= xLDY;
  default_le <= eZERO;
  admode <= sEINDIRECT;
when "0110100001" =>          -- $a1, LEA Zeropage indexed with X indirect 16bit: (zp,X)  (65k)
  operation <= xLEA;
  idxreg <= iXR;
  indwidth <= wWORD;
  parwidth <= pBYTE;
  admode <= sPREINDIRECT;
when "0110100010" =>          -- $a2, LDX E indirect: (E)  (65k)
  operation <= xLDX;
  default_le <= eZERO;
  admode <= sEINDIRECT;
when "0110100100" =>          -- $a4, INV Accumulator:   (65k)
  operation <= xINV_A;
  admode <= sIMPLIED;
when "0110100101" =>          -- $a5, SBE Immediate: #byte  (65k)
  operation <= xSBE;
  parwidth <= pw_rs;
  admode <= sIMMEDIATE;
when "0110101000" =>          -- $a8, SAB Implied:   (65k)
  operation <= xSAB;
  admode <= sIMPLIED;
when "0110101001" =>          -- $a9, LDA E indirect: (E)  (65k)
  operation <= xLDA;
  default_le <= eZERO;
  admode <= sEINDIRECT;
when "0110101101" =>          -- $ad, PEA Absolute 16bit: abs  (65k)
  operation <= xPEA;
  parwidth <= pw_wq;
  admode <= sABSOLUTE;
when "0110101110" =>          -- $ae, LEA Absolute 16bit: abs  (65k)
  operation <= xLEA;
  parwidth <= pw_wq;
  admode <= sABSOLUTE;
when "0110110001" =>          -- $b1, LEA Zeropage indirect 16bit indexed with Y: (zp),Y  (65k)
  operation <= xLEA;
  idxreg <= iYR;
  indwidth <= wWORD;
  parwidth <= pBYTE;
  admode <= sPOSTINDIRECT;
when "0110110010" =>          -- $b2, LEA Zeropage indirect 16bit: (zp)  (65k)
  operation <= xLEA;
  indwidth <= wWORD;
  parwidth <= pBYTE;
  admode <= sINDIRECT;
when "0110110100" =>          -- $b4, BCN Accumulator:   (65k)
  operation <= xBCN_A;
  admode <= sIMPLIED;
when "0110110101" =>          -- $b5, SBE Accumulator:   (65k)
  operation <= xSBE_A;
  admode <= sIMPLIED;
when "0110111000" =>          -- $b8, SEB Implied:   (65k)
  operation <= xSEB;
  admode <= sIMPLIED;
when "0110111001" =>          -- $b9, LEA Absolute 16bit indexed with Y: abs,Y  (65k)
  operation <= xLEA;
  idxreg <= iYR;
  parwidth <= pw_wq;
  admode <= sABSOLUTEIND;
when "0110111010" =>          -- $ba, SAX Implied:   (65k)
  operation <= xSAX;
  admode <= sIMPLIED;
when "0110111101" =>          -- $bd, PEA Absolute 16bit indexed with X: abs,X  (65k)
  operation <= xPEA;
  idxreg <= iXR;
  parwidth <= pw_wq;
  admode <= sABSOLUTEIND;
when "0110111110" =>          -- $be, LEA Absolute 16bit indexed with X: abs,X  (65k)
  operation <= xLEA;
  idxreg <= iXR;
  parwidth <= pw_wq;
  admode <= sABSOLUTEIND;
when "0111000000" =>          -- $c0, CPY E indirect: (E)  (65k)
  operation <= xCPY;
  admode <= sEINDIRECT;
when "0111000010" =>          -- $c2, PEA Absolute indirect 16bit indexed with Y: (abs),Y  (65k)
  operation <= xPEA;
  idxreg <= iYR;
  indwidth <= wWORD;
  parwidth <= pWORD;
  admode <= sPOSTINDIRECT;
when "0111000100" =>          -- $c4, EXT Accumulator:   (65k)
  operation <= xEXT_A;
  admode <= sIMPLIED;
when "0111000101" =>          -- $c5, SBS Immediate: #byte  (65k)
  operation <= xSBS;
  parwidth <= pw_rs;
  admode <= sIMMEDIATE;
when "0111001000" =>          -- $c8, TPA Implied:   (65k)
  operation <= xTPA;
  admode <= sIMPLIED;
when "0111001001" =>          -- $c9, CMP E indirect: (E)  (65k)
  operation <= xCMP;
  admode <= sEINDIRECT;
when "0111001010" =>          -- $ca, TSY Implied:   (65k)
  operation <= xTSY;
  admode <= sIMPLIED;
when "0111001101" =>          -- $cd, DEC E indirect: (E)  (65k)
  operation <= xDEC;
  admode <= sEINDIRECT;
when "0111010100" =>          -- $d4, SWP Accumulator:   (65k)
  operation <= xSWP_A;
  admode <= sIMPLIED;
when "0111010101" =>          -- $d5, SBS Accumulator:   (65k)
  operation <= xSBS_A;
  admode <= sIMPLIED;
when "0111011000" =>          -- $d8, SAE Implied:   (65k)
  operation <= xSAE;
  admode <= sIMPLIED;
when "0111011010" =>          -- $da, SAY Implied:   (65k)
  operation <= xSAY;
  admode <= sIMPLIED;
when "0111011100" =>          -- $dc, JSR Address Long: long 
  operation <= xJSR;
  default_le <= eSIGN;
  parwidth <= pLONG;
  admode <= sADDR;
when "0111100000" =>          -- $e0, CPX E indirect: (E)  (65k)
  operation <= xCPX;
  admode <= sEINDIRECT;
when "0111100010" =>          -- $e2, PEA Absolute indexed with X indirect 16bit: (abs,X)  (65k)
  operation <= xPEA;
  idxreg <= iXR;
  indwidth <= wWORD;
  parwidth <= pWORD;
  admode <= sPREINDIRECT;
when "0111100100" =>          -- $e4, RMB E indirect: (E)  (65k)
  operation <= xRMB;
  admode <= sEINDIRECT;
when "0111100101" =>          -- $e5, SBB Immediate: #byte  (65k)
  operation <= xSBB;
  parwidth <= pw_rs;
  admode <= sIMMEDIATE;
when "0111101000" =>          -- $e8, TAB Implied:   (65k)
  operation <= xTAB;
  admode <= sIMPLIED;
when "0111101001" =>          -- $e9, SBC E indirect: (E)  (65k)
  operation <= xSBC;
  admode <= sEINDIRECT;
when "0111101010" =>          -- $ea, TEB Implied:   (65k)
  operation <= xTEB;
  admode <= sIMPLIED;
when "0111101101" =>          -- $ed, INC E indirect: (E)  (65k)
  operation <= xINC;
  admode <= sEINDIRECT;
when "0111110100" =>          -- $f4, WMB E indirect: (E)  (65k)
  operation <= xWMB;
  admode <= sEINDIRECT;
when "0111110101" =>          -- $f5, SBB Accumulator:   (65k)
  operation <= xSBB_A;
  admode <= sIMPLIED;
when "0111111000" =>          -- $f8, TBA Implied:   (65k)
  operation <= xTBA;
  admode <= sIMPLIED;
when "0111111010" =>          -- $fa, TBE Implied:   (65k)
  operation <= xTBE;
  admode <= sIMPLIED;
when others =>
  is_valid <= '0';
end case;

end process;

end Behavioral;

